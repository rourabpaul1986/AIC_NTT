

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Helper utility package: clog2 and simple helpers
package util_pkg is
  -- ceiling(log2) for natural > 0
  function clog2(n : natural) return natural;
end package util_pkg;

package body util_pkg is
  function clog2(n : natural) return natural is
    variable v : natural := n - 1;
    variable c : natural := 0;
  begin
    if n <= 1 then
      return 1;
    end if;
    while v > 0 loop
      v := v / 2;
      c := c + 1;
    end loop;
    return c;
  end function clog2;
end package body util_pkg;

use work.util_pkg.all;

-- Main entity
entity NTTCore is
  generic (
    -- Top-level configuration (kept similar to original SV generics)
    NTT            : natural := 1;
    LOGQ           : natural := 28;
    LOGN           : natural := 11;
    PE             : natural := 8;

    NTT_TYPE       : string  := "mfntt_dit_nr-mintt_dif_rn";
    Q_VALUE        : natural := 0;
    WORD_SIZE      : natural := 12;

    ADD_LAT        : natural := 1;
    INTMUL_LAT     : natural := 2;
    INTMUL_TYPE    : string  := "fpga_dsp";
    MODRED_TYPE    : string  := "default";
    MODRED_LAT     : natural := 1;
    MODRED_COREMUL_LAT : natural := 1;

    INSTANTIATE_MULT_ADD : natural := 0;
    NUM_POLY_MEMS  : natural := 1;

    MEMORY_OPTIMIZED : natural := 0;
    TW_ROM_MEM_TYPE : string := "fpga_block";
    ROM_ADDR_WIDTH  : natural := 32;
    RAM_RD_LAT      : natural := 2;
    ROM_RD_LAT      : natural := 2;

    NO_BFU         : natural := 0;


    ADDR_WIDTH     : natural := clog2((NUM_POLY_MEMS * (2 ** LOGN)) / 2 / PE)
  );
  port (
    clk      : in  std_logic;
    rst      : in  std_logic;
    forward  : in  std_logic;
    opcode   : in  std_logic_vector(1 downto 0);

    q                : in  std_logic_vector(LOGQ-1 downto 0);
    montgomery_factor: in  std_logic_vector(LOGQ-1 downto 0);
    rom_base_addr    : in  std_logic_vector(ROM_ADDR_WIDTH-1 downto 0);

    ram_wen  : out std_logic;
    ram_raddr: out std_logic_vector(ADDR_WIDTH-1 downto 0);
    ram_waddr: out std_logic_vector(ADDR_WIDTH-1 downto 0);

    -- flattened ram read data: layout: for g in 0..PE-1, for pair in 0..1
    -- bit-width = PE * 2 * LOGQ
    ram_rdata_flat : in  std_logic_vector((PE*2*LOGQ)-1 downto 0);
    ram_wdata_flat : out std_logic_vector((PE*2*LOGQ)-1 downto 0);

    poly_base_a : in  std_logic_vector(util_pkg.clog2(NUM_POLY_MEMS)-1 downto 0);
    poly_base_b : in  std_logic_vector(util_pkg.clog2(NUM_POLY_MEMS)-1 downto 0);

    done : out std_logic
  );
end entity NTTCore;

architecture rtl of NTTCore is
  -- conveniences:
  subtype word_t is std_logic_vector(LOGQ-1 downto 0);
  constant N : natural := 2 ** LOGN;

  -- Internal signals (mirroring SV names)
  signal rom_base_addr_reg : std_logic_vector(ROM_ADDR_WIDTH-1 downto 0);
  signal forward_internal  : std_logic;

  -- Control/status
  signal ntt_opcode, add_opcode, sub_opcode, mult_opcode : std_logic;
  signal montgomery_factor_DP : std_logic_vector(LOGQ-1 downto 0);
  signal poly_base_a_DP, poly_base_b_DP : std_logic_vector(util_pkg.clog2(NUM_POLY_MEMS)-1 downto 0);

  -- Address generation and control signals (many of these are placeholders)
  signal rst_addr_gen_nr, rst_addr_gen_rn : std_logic;
  signal done_nr, done_rn, done_internal, done_polyArith : std_logic;
  signal ident_store_nr, ident_store_rn, ident_store : std_logic;
  signal ident_store_delayed : std_logic;
  signal rd_addr_nr, rd_addr_rn, rd_addr, rd_addr_delayed : std_logic_vector(ADDR_WIDTH-1 downto 0);
  signal dest_rom_gap_nr, dest_rom_gap_rn, dest_rom_gap, dest_rom_gap_delayed : std_logic_vector(util_pkg.clog2(PE) downto 0);

  -- Poly arith block signals
  signal raddr_polyArith : std_logic_vector((util_pkg.clog2(NUM_POLY_MEMS)+ADDR_WIDTH)-1 downto 0);
  signal waddr_polyArith : std_logic_vector((util_pkg.clog2(NUM_POLY_MEMS)+ADDR_WIDTH)-1 downto 0);
  signal bf_a_polyArith_flat : std_logic_vector((PE*LOGQ)-1 downto 0);
  signal bf_b_polyArith_flat : std_logic_vector((PE*LOGQ)-1 downto 0);
  signal bf_c_polyArith_flat : std_logic_vector((PE*LOGQ)-1 downto 0);
  signal dest_rom_gap_PolyArith : std_logic_vector(util_pkg.clog2(PE) downto 0);
  signal ident_store_PolyArith, swap_store_PolyArith, valid_PolyArith : std_logic;

  -- Twiddle factor outputs (flattened)
  signal tw_flat : std_logic_vector((PE*LOGQ)-1 downto 0);

  -- Butterfly outputs flattened: for each PE, two words
  signal btf_out_flat : std_logic_vector((PE*2*LOGQ)-1 downto 0);

  -- store signals
  signal valid_delayed : std_logic;
  signal wen : std_logic;
  signal waddr : std_logic_vector(ADDR_WIDTH-1 downto 0);
  signal wdata_flat : std_logic_vector((PE*2*LOGQ)-1 downto 0);

  -- done DP flag
  signal done_DP : std_logic := '0';

  -- temporary control
  signal done_tmp : std_logic;

  -- helper functions to index flattened vectors
  impure function idx_word_flat(flat : std_logic_vector; i : natural) return std_logic_vector is
    variable start_bit : integer := flat'left - integer(i)*integer(LOGQ);
    variable res : std_logic_vector(LOGQ-1 downto 0);
  begin
    res := flat(start_bit downto start_bit - integer(LOGQ) + 1);
    return res;
  end function idx_word_flat;


begin


  process(clk)
  begin
    if rising_edge(clk) then
      rom_base_addr_reg <= rom_base_addr;
    end if;
  end process;


  process(clk)
  begin
    if rising_edge(clk) then
      forward_internal <= forward;
    end if;
  end process;

  -- Input registers and op selection (registered on clk)
  process(clk)
  begin
    if rising_edge(clk) then
      poly_base_a_DP <= poly_base_a;
      poly_base_b_DP <= poly_base_b;
      montgomery_factor_DP <= montgomery_factor;
      -- ntt_opcode and arithmetic op decode:
      if INSTANTIATE_MULT_ADD = 0 then
        ntt_opcode <= '1'; -- only NTT
      else
        -- when INSTANTIATE_MULT_ADD = 1, opcode values decide
        ntt_opcode <= (opcode = "00") ? '1' : '0'; -- emulate: opcode==0 => NTT
      end if;
      mult_opcode <= (INSTANTIATE_MULT_ADD /= 0 and opcode = "01") ? '1' : '0';
      add_opcode  <= (INSTANTIATE_MULT_ADD /= 0 and opcode = "10") ? '1' : '0';
      sub_opcode  <= (INSTANTIATE_MULT_ADD /= 0 and opcode = "11") ? '1' : '0';
    end if;
  end process;

  --------------------------------------------------------------------

  --------------------------------------------------------------------
  component AddrGen
    generic (
      LOGN_g : natural;
      PE_g   : natural;
      LATENCY_g : natural;
      IS_NR_g  : natural
    );
    port (
      clk  : in  std_logic;
      rst  : in  std_logic;
      ident_store : in std_logic;
      dest_rom_gap : in std_logic_vector(util_pkg.clog2(PE) downto 0);
      done : out std_logic;
      addr_out : out std_logic_vector(ADDR_WIDTH-1 downto 0)
    );
  end component;

  component AddrGen_PolyArith
    generic (
      LOGN_g : natural;
      PE_g   : natural;
      BTF_TYPE_g : string;
      NUM_POLY_g : natural;
      BFU_LAT_g : natural;
      SHUFFLER_LAT_g : natural;
      BRAM_RD_LAT_g : natural
    );
    port (
      clk  : in std_logic;
      rst  : in std_logic;
      sub_opcode : in std_logic;
      poly_base_a : in std_logic_vector((util_pkg.clog2(NUM_POLY_MEMS)+ADDR_WIDTH)-1 downto 0);
      poly_base_b : in std_logic_vector((util_pkg.clog2(NUM_POLY_MEMS)+ADDR_WIDTH)-1 downto 0);
      valid : out std_logic;
      swap  : out std_logic;
      done  : out std_logic;
      addr_out : out std_logic_vector((util_pkg.clog2(NUM_POLY_MEMS)+ADDR_WIDTH)-1 downto 0)
    );
  end component;

  component DataShuffler_PolyArith
    generic (
      BTF_TYPE_g : string;
      LOGN_g : natural;
      LOGQ_g : natural;
      PE_g   : natural;
      NUM_POLY_g : natural;
      BRAM_RD_LAT_g : natural;
      ADD_SUB_LAT_g : natural;
      BFU_LAT_g : natural
    );
    port (
      clk  : in std_logic;
      rst  : in std_logic;
      opcode : in std_logic_vector(1 downto 0);
      valid_in : in std_logic;
      montgomery_factor : in std_logic_vector(LOGQ-1 downto 0);
      swap : in std_logic;
      addr : in std_logic_vector((util_pkg.clog2(NUM_POLY_MEMS)+ADDR_WIDTH)-1 downto 0);
      rdata_flat : in std_logic_vector((PE*2*LOGQ)-1 downto 0);
      bf_a_flat : out std_logic_vector((PE*LOGQ)-1 downto 0);
      bf_b_flat : out std_logic_vector((PE*LOGQ)-1 downto 0);
      bf_c_flat : out std_logic_vector((PE*LOGQ)-1 downto 0);
      ident_store : out std_logic;
      swap_store  : out std_logic;
      dest_rom_gap : out std_logic_vector(util_pkg.clog2(PE) downto 0);
      waddr : out std_logic_vector((util_pkg.clog2(NUM_POLY_MEMS)+ADDR_WIDTH)-1 downto 0);
      valid_out : out std_logic
    );
  end component;

  component TwiddleGen
    generic (
      NTT_g : natural;
      LOGQ_g : natural;
      LOGN_g : natural;
      PE_g : natural;
      MEMORY_OPTIMIZED_g : natural;
      NTT_TYPE_g : string;
      ROM_RD_LAT_g : natural;
      ROM_ADDR_WIDTH_g : natural;
      MEM_TYPE_g : string;
      INTMUL_LAT_g : natural;
      INTMUL_TYPE_g : string;
      Q_VALUE_g : natural;
      WORD_SIZE_g : natural;
      MODRED_LAT_g : natural;
      MODRED_TYPE_g : string;
      MODRED_L_g : natural;
      MODRED_COREMUL_LAT_g : natural
    );
    port (
      clk  : in std_logic;
      rst  : in std_logic;
      forward : in std_logic;
      rom_base_addr : in std_logic_vector(ROM_ADDR_WIDTH-1 downto 0);
      q : in std_logic_vector(LOGQ-1 downto 0);
      tw_out_flat : out std_logic_vector((PE*LOGQ)-1 downto 0)
    );
  end component;

  component shiftreg
    generic (
      DELAY_g : natural;
      LOGQ_g  : natural
    );
    port (
      clk : in std_logic;
      data_in : in std_logic_vector(LOGQ_g-1 downto 0);
      data_out: out std_logic_vector(LOGQ_g-1 downto 0)
    );
  end component;

  component btf_uni
    generic (
      LOGQ_g : natural;
      Q_VALUE_g : natural;
      WORD_SIZE_g : natural;
      MODADD_LAT_g : natural;
      INTMUL_LAT_g : natural;
      INTMUL_TYPE_g : string;
      MODRED_LAT_g : natural;
      MODRED_TYPE_g : string;
      MODRED_L_g : natural;
      MODRED_COREMUL_LAT_g : natural;
      BTF_TYPE_g : string;
      SHIFT_AE_g : natural;
      DIV_BY_2_g : natural
    );
    port (
      clk : in std_logic;
      dif_dit : in std_logic;
      div_by_2 : in std_logic;
      opcode : in std_logic_vector(1 downto 0);
      q : in std_logic_vector(LOGQ_g-1 downto 0);
      a : in std_logic_vector(LOGQ_g-1 downto 0);
      b : in std_logic_vector(LOGQ_g-1 downto 0);
      w : in std_logic_vector(LOGQ_g-1 downto 0);
      e : out std_logic_vector(LOGQ_g-1 downto 0);
      o : out std_logic_vector(LOGQ_g-1 downto 0)
    );
  end component;

  component FFTButterfly
    generic (
      BTF_TYPE_g : string;
      DIV_BY_2_g : natural
    );
    port (
      clk : in std_logic;
      dif_dit : in std_logic;
      div_by_2 : in std_logic;
      opcode : in std_logic_vector(1 downto 0);
      a : in std_logic_vector(LOGQ-1 downto 0);
      b : in std_logic_vector(LOGQ-1 downto 0);
      w : in std_logic_vector(LOGQ-1 downto 0);
      e : out std_logic_vector(LOGQ-1 downto 0);
      o : out std_logic_vector(LOGQ-1 downto 0)
    );
  end component;

  component DataShuffler
    generic (
      LOGQ_g : natural;
      LOGN_g : natural;
      PE_g : natural
    );
    port (
      clk  : in std_logic;
      valid : in std_logic;
      ident_store : in std_logic;
      dest_rom_gap : in std_logic_vector(util_pkg.clog2(PE) downto 0);
      swap_store : in std_logic;
      is_poly_arith : in std_logic;
      bf_rd_addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
      bf_data_flat : in std_logic_vector((PE*2*LOGQ)-1 downto 0);
      wen : out std_logic;
      waddr : out std_logic_vector(ADDR_WIDTH-1 downto 0);
      wdata_flat : out std_logic_vector((PE*2*LOGQ)-1 downto 0)
    );
  end component;

  --------------------------------------------------------------------
  -- Instantiations: address generators, twiddle gen, data shufflers, BF units
  --------------------------------------------------------------------

  -- AddrGen instances (NR and RN) when needed:
  addr_gen_nr_inst : if true generate
    -- instantiate only if NR path exists in higher-level design
    begin
      AG_NR: AddrGen
       generic map (
         LOGN_g => LOGN,
         PE_g => PE,
         LATENCY_g => 1,
         IS_NR_g => 1
       )
       port map (
         clk => clk,
         rst => rst_addr_gen_nr,
         ident_store => ident_store_nr,
         dest_rom_gap => dest_rom_gap_nr,
         done => done_nr,
         addr_out => rd_addr_nr
       );
  end generate;

  addr_gen_rn_inst : if true generate
    AG_RN: AddrGen
       generic map (
         LOGN_g => LOGN,
         PE_g => PE,
         LATENCY_g => 1,
         IS_NR_g => 0
       )
       port map (
         clk => clk,
         rst => rst_addr_gen_rn,
         ident_store => ident_store_rn,
         dest_rom_gap => dest_rom_gap_rn,
         done => done_rn,
         addr_out => rd_addr_rn
       );
  end generate;

  -- Twiddle generator:
  tw_gen_inst : TwiddleGen
    generic map (
      NTT_g => NTT,
      LOGQ_g => LOGQ,
      LOGN_g => LOGN,
      PE_g => PE,
      MEMORY_OPTIMIZED_g => MEMORY_OPTIMIZED,
      NTT_TYPE_g => NTT_TYPE,
      ROM_RD_LAT_g => ROM_RD_LAT,
      ROM_ADDR_WIDTH_g => ROM_ADDR_WIDTH,
      MEM_TYPE_g => TW_ROM_MEM_TYPE,
      INTMUL_LAT_g => INTMUL_LAT,
      INTMUL_TYPE_g => INTMUL_TYPE,
      Q_VALUE_g => Q_VALUE,
      WORD_SIZE_g => WORD_SIZE,
      MODRED_LAT_g => MODRED_LAT,
      MODRED_TYPE_g => MODRED_TYPE,
      MODRED_L_g => natural( (LOGQ + WORD_SIZE - 1) / WORD_SIZE ),
      MODRED_COREMUL_LAT_g => MODRED_COREMUL_LAT
    )
    port map (
      clk => clk,
      rst => rst_addr_gen_nr, -- tie to a reset; adjust per timing logic
      forward => forward_internal,
      rom_base_addr => rom_base_addr_reg,
      q => q,
      tw_out_flat => tw_flat
    );

  -- Butterfly instantiation loop
  gen_bfs : for g in 0 to PE-1 generate
    -- Extract per-PE inputs from flattened ram_rdata or poly arith outputs
    signal a_in, b_in, w_in : std_logic_vector(LOGQ-1 downto 0);
    signal e_out, o_out : std_logic_vector(LOGQ-1 downto 0);
  begin
    -- Extract read operands for this PE when NTT path: we assume ram_rdata_flat
    a_in <= ram_rdata_flat((PE*2*LOGQ)-1 - (g*2*LOGQ) downto (PE*2*LOGQ) - (g*2*LOGQ) - LOGQ + 1)
             when ntt_opcode = '1' else bf_a_polyArith_flat((g+1)*LOGQ-1 downto g*LOGQ);
    b_in <= ram_rdata_flat((PE*2*LOGQ)-1 - (g*2*LOGQ + LOGQ) downto (PE*2*LOGQ) - (g*2*LOGQ + LOGQ) - LOGQ + 1)
             when ntt_opcode = '1' else bf_b_polyArith_flat((g+1)*LOGQ-1 downto g*LOGQ);
    w_in <= tw_flat((g+1)*LOGQ-1 downto g*LOGQ) when ntt_opcode = '1' else bf_c_polyArith_flat((g+1)*LOGQ-1 downto g*LOGQ);

    -- Choose BF implementation: btf_uni (NTT) or FFTButterfly (FFT)
    btf_inst : if NO_BFU = 0 generate
      btf_u : btf_uni
        generic map (
          LOGQ_g => LOGQ,
          Q_VALUE_g => Q_VALUE,
          WORD_SIZE_g => WORD_SIZE,
          MODADD_LAT_g => ADD_LAT,
          INTMUL_LAT_g => INTMUL_LAT,
          INTMUL_TYPE_g => INTMUL_TYPE,
          MODRED_LAT_g => MODRED_LAT,
          MODRED_TYPE_g => MODRED_TYPE,
          MODRED_L_g => natural((LOGQ + WORD_SIZE - 1) / WORD_SIZE),
          MODRED_COREMUL_LAT_g => MODRED_COREMUL_LAT,
          BTF_TYPE_g => "unified",
          SHIFT_AE_g => 1,
          DIV_BY_2_g => (IS_INVERSE or (NTT_TYPE = "mfntt_dit_nr-mintt_dif_rn")) ? 1 : 0
        )
        port map (
          clk => clk,
          dif_dit => '0', -- do_dit derivation omitted for brevity
          div_by_2 => '0',
          opcode => opcode,
          q => q,
          a => a_in,
          b => b_in,
          w => w_in,
          e => e_out,
          o => o_out
        );
    end generate;

    -- For NO_BFU = 1 a simple shift-through (delay) could be instantiated; omitted.

    -- Pack outputs back into the flat btf_out_flat
    -- We place `e_out` and `o_out` at positions corresponding to `g`
    btf_out_flat((g*2+1)*LOGQ-1 downto (g*2)*LOGQ) <= e_out & o_out; -- note: pack may require reorder
  end generate;

  -- Address/valid delay registers and data shuffler
  -- Simplified: we directly call DataShuffler, and tie valid/waddr/wdata outputs
  data_shuffler_inst : DataShuffler
    generic map (
      LOGQ_g => LOGQ,
      LOGN_g => LOGN,
      PE_g => PE
    )
    port map (
      clk => clk,
      valid => valid_delayed,
      ident_store => ident_store_delayed,
      dest_rom_gap => dest_rom_gap_delayed,
      swap_store => swap_store_PolyArith,
      is_poly_arith => (ntt_opcode = '0'),
      bf_rd_addr => rd_addr_delayed,
      bf_data_flat => btf_out_flat,
      wen => wen,
      waddr => waddr,
      wdata_flat => wdata_flat
    );

  -- Connect the flattened wdata to external ram_wdata_flat (gated by wen and done_DP)
  ram_wdata_flat <= wdata_flat;
  ram_wen <= wen and not done_DP;

  -- ram raddr/waddr logic (simplified)
  ram_raddr <= rd_addr; -- drive directly; in original this depends on NUM_POLY_MEMS etc.
  ram_waddr <= waddr;

  -- done signalling: delayed version of done_internal
  done_tmp <= done_internal; -- ideally this is delayed by BTF_LAT+RAM_RD_LAT+... but omitted here
  done <= done_tmp;

  -- done_DP register
  process(clk)
  begin
    if rising_edge(clk) then
      if rst = '1' then
        done_DP <= '0';
      elsif done = '1' then
        done_DP <= '1';
      end if;
    end if;
  end process;



end architecture rtl;
